--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x:2
-- 	 network size y:2
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.TB_Package.all;

USE ieee.numeric_std.ALL;
--use IEEE.math_real."ceil";
--use IEEE.math_real."log2";

entity tb_network_2x2 is
port(
    clk : in std_logic;
    reset : in std_logic;
    uart_read_0 : in std_logic;
    uart_read_1 : in std_logic;
    uart_read_2 : in std_logic;
    uart_read_3 : in std_logic;
    uart_write_0 : out std_logic;
    uart_write_1 : out std_logic;
    uart_write_2 : out std_logic;
    uart_write_3 : out std_logic;
    TX_L_0_out: out std_logic_vector(31 downto 0);
    TX_L_1_out: out std_logic_vector(31 downto 0);
    TX_L_2_out: out std_logic_vector(31 downto 0);
    TX_L_3_out: out std_logic_vector(31 downto 0)
   );
end tb_network_2x2;


architecture behavior of tb_network_2x2 is

-- Declaring network component
component network_2x2 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic;
	clk: in  std_logic;
	Rxy_reconf: in  std_logic_vector(7 downto 0);
	Reconfig : in std_logic;
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0)

            );
end component;
component NoC_Node is
generic( current_address : integer := 0; stim_file: string :="code.txt");
port( reset        : in std_logic;
      clk          : in std_logic;
      uart_read : in std_logic;
      uart_write : out std_logic;

        credit_in : in std_logic;
        valid_out: out std_logic;
        TX: out std_logic_vector(31 downto 0);

        credit_out : out std_logic;
        valid_in: in std_logic;
        RX: in std_logic_vector(31 downto 0)
   );
end component; --component NoC_Node

-- generating bulk signals...
	signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
	signal credit_counter_out_0:  std_logic_vector (1 downto 0);
	signal credit_out_L_0, credit_in_L_0, valid_in_L_0, valid_out_L_0: std_logic;
	signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
	signal credit_counter_out_1:  std_logic_vector (1 downto 0);
	signal credit_out_L_1, credit_in_L_1, valid_in_L_1, valid_out_L_1: std_logic;
	signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
	signal credit_counter_out_2:  std_logic_vector (1 downto 0);
	signal credit_out_L_2, credit_in_L_2, valid_in_L_2, valid_out_L_2: std_logic;
	signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
	signal credit_counter_out_3:  std_logic_vector (1 downto 0);
	signal credit_out_L_3, credit_in_L_3, valid_in_L_3, valid_out_L_3: std_logic;
	--------------

signal Rxy_reconf: std_logic_vector (7 downto 0) := "01111101";
signal Reconfig: std_logic := '0';
 constant clk_period : time := 1 ns;
signal not_reset : std_logic :='0';

-- Those are going out. later I will multiplex them, so that all of them will be able to communicate with physical uart.
 -- signal uart_read_0   : std_logic;
 -- signal uart_read_1   : std_logic;
 -- signal uart_read_2   : std_logic;
 -- signal uart_read_3   : std_logic;
 --
 -- signal uart_write_0  : std_logic;
 -- signal uart_write_1  : std_logic;
 -- signal uart_write_2  : std_logic;
 -- signal uart_write_3  : std_logic;

begin
TX_L_0_out <=TX_L_0;
TX_L_1_out <=TX_L_1;
TX_L_2_out <=TX_L_2;
TX_L_3_out <=TX_L_3;
-- instantiating the network
NoC: network_2x2 generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk, Rxy_reconf, Reconfig,
	--------------
	RX_L_0, credit_out_L_0, valid_out_L_0, credit_in_L_0, valid_in_L_0,  TX_L_0,
	--------------
	RX_L_1, credit_out_L_1, valid_out_L_1, credit_in_L_1, valid_in_L_1,  TX_L_1,
	--------------
	RX_L_2, credit_out_L_2, valid_out_L_2, credit_in_L_2, valid_in_L_2,  TX_L_2,
	--------------
	RX_L_3, credit_out_L_3, valid_out_L_3, credit_in_L_3, valid_in_L_3,  TX_L_3
            );
not_reset <= not reset;

-- connecting the PEs
PE_0: NoC_Node
generic map( current_address => 0, stim_file => "/home/tsotnep/ownCloud/git/Bonfire/tmp/simul_temp/code_0.txt")
port map( not_reset, clk,
uart_read => uart_read_0,
uart_write => uart_write_0,

        credit_in => credit_out_L_0,
        valid_out => valid_in_L_0,
        TX => RX_L_0,

        credit_out => credit_in_L_0,
        valid_in => valid_out_L_0,
        RX => TX_L_0
   );
PE_1: NoC_Node
generic map( current_address => 1, stim_file => "/home/tsotnep/ownCloud/git/Bonfire/tmp/simul_temp/code_1.txt")
port map( not_reset, clk,
uart_read => uart_read_1,
uart_write => uart_write_1,

        credit_in => credit_out_L_1,
        valid_out => valid_in_L_1,
        TX => RX_L_1,

        credit_out => credit_in_L_1,
        valid_in => valid_out_L_1,
        RX => TX_L_1
   );
PE_2: NoC_Node
generic map( current_address => 2, stim_file => "/home/tsotnep/ownCloud/git/Bonfire/tmp/simul_temp/code_2.txt")
port map( not_reset, clk,
uart_read => uart_read_2,
uart_write => uart_write_2,

        credit_in => credit_out_L_2,
        valid_out => valid_in_L_2,
        TX => RX_L_2,

        credit_out => credit_in_L_2,
        valid_in => valid_out_L_2,
        RX => TX_L_2
   );
PE_3: NoC_Node
generic map( current_address => 3, stim_file => "/home/tsotnep/ownCloud/git/Bonfire/tmp/simul_temp/code_3.txt")
port map( not_reset, clk,
uart_read => uart_read_3,
uart_write => uart_write_3,

        credit_in => credit_out_L_3,
        valid_out => valid_in_L_3,
        TX => RX_L_3,

        credit_out => credit_in_L_3,
        valid_in => valid_out_L_3,
        RX => TX_L_3
   );



end;
